module MutEx #(parameter N)(
  input  ipClk,
  input  ipReset,

  input  [N-1:0]ipRequest,
  output [N-1:0]opGrant
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

