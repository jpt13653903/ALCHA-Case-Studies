module ADS7056(
  input        ipClk,
  input        ipReset,

  output       opSClk,
  output       opnCS,
  input        ipData,

  output [13:0]opData,
  output       opValid
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

