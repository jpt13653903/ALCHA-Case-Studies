module MasterTriggerGen(
  input  ipClk,
  input  ipReset,

  input  ipPeriod,
  output opTrigger
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

