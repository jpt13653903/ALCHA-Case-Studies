module PlaceHolder(
  input ipClk,
  input ipReset
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

