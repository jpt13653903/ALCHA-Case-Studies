module RealWindow(
  input  ipClk,
  input  ipReset,

  input  PACKET ipInput,
  output opReady,

  output DATA_PACKET opOutput,
  input  ipReady
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

