module TriggerDelay(
  input       ipClk,
  input       ipReset,

  input       ipEnable,
  input [31:0]ipDelay,
  input [31:0]ipLength,

  input       ipTrigger,
  output      opTrigger
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

