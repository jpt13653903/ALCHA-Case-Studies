module IQ_Window(
  input  ipClk,
  input  ipReset,

  input  IQ_PACKET ipInput,
  output opReady,

  output IQ_PACKET opOutput,
  input  ipReady
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

