module RealFFT(
  input  ipClk,
  input  ipReset,

  input  DATA_PACKET ipInput,
  output opReady,

  output IQ_PACKET opOutput,
  input  ipReady
);
//------------------------------------------------------------------------------

endmodule
//------------------------------------------------------------------------------

